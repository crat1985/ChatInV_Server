module utils

import db.sqlite

pub fn ask_credentials(mut user &User, db sqlite.DB) (string, string, string) {
	for {
		mut data := []u8{len: 1024}
		user.write_string("Pseudo : ") or {
			return "Error while asking pseudo : $err", "", ""
		}
		mut lenght := user.read(mut data) or {
			return "Error while reading pseudo : $err", "", ""
		}
		mut pseudo := data[0..lenght].bytestr()
		user.write_string("Password : ") or {
			return "Error while asking password : $err", "", ""
		}
		data = []u8{len: 1024}
		lenght = user.read(mut data) or {
			return "Error while reading password : $err", "", ""
		}
		mut password := data[0..lenght].bytestr()
		if pseudo.len < 8 || password.len < 8 {
			println("[LOG] ${user.peer_ip() or {"IPERROR"}} => 'Pseudo or password too short !'")
			user.write_string("Pseudo or password too short !\n") or {
				return "Error while writing too short error : $err", "", ""
			}
			continue
		}

		account := get_account_by_pseudo(db, pseudo)
		if password == account.password {
			return "", pseudo, password
		}

		println("[LOG] ${user.peer_ip() or {"IPERROR"}} => 'Wrong password !'")
		user.write_string("Wrong password !\n") or {
			return "Error while sending 'Wrong password' to ${user.peer_ip() or {"IPERROR"}}", "", ""
		}
	}

	return "This could never happens !", "", ""

}
